`timescale 1ns/1ns
`include "lab3A.v"
module lab3A_tb(); 
reg A,B,C,D;
wire f;
lab3A ab(A,B,C,D,f);
initial
begin
$dumpfile("lab3A_tb.vcd");
$dumpvars(0, lab3A_tb);
A=1'b0; B=1'b0; C=1'b0; D=1'b0;
#20;
A=1'b0;B=1'b0;C=1'b0;D=1'b1;
#20;
A=1'b0;B=1'b0;C=1'b1;D=1'b0;
#20;
A=1'b0;B=1'b0;C=1'b1;D=1'b1;
#20;
A=1'b0;B=1'b1;C=1'b0;D=1'b0;
#20;
A=1'b0;B=1'b1;C=1'b0;D=1'b1;
#20;
A=1'b0;B=1'b1;C=1'b1;D=1'b0;
#20;
A=1'b0;B=1'b1;C=1'b1;D=1'b1;
#20;
A=1'b1;B=1'b0;C=1'b0;D=1'b0;
#20;
A=1'b1;B=1'b0;C=1'b0;D=1'b1;
#20;
A=1'b1;B=1'b0;C=1'b1;D=1'b0;
#20;
A=1'b1;B=1'b0;C=1'b1;D=1'b1;
#20;
A=1'b1;B=1'b1;C=1'b0;D=1'b0;
#20;
A=1'b0;B=1'b1;C=1'b0;D=1'b1;
#20;
A=1'b1;B=1'b1;C=1'b1;D=1'b0;
#20;
A=1'b1;B=1'b1;C=1'b1;D=1'b1;
#20;
$display("Test Complete");
end
endmodule
